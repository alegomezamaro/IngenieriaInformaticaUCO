** Profile: "SCHEMATIC1-S4"  [ C:\Users\gomez\Desktop\S4\S4-PSpiceFiles\SCHEMATIC1\S4.sim ] 

** Creating circuit file "S4.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.STMLIB "../../../s4-pspicefiles/s4.stl" 
* From [PSPICE NETLIST] section of C:\Users\gomez\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 3200ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
